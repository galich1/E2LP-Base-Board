--------------------------------------------------------------------------------
-- Company: 
-- Engineer:
--
-- Create Date:   12:00:15 03/19/2021
-- Design Name:   
-- Module Name:   C:/LRI2/UartController/UARTtb.vhd
-- Project Name:  UartController
-- Target Device:  
-- Tool versions:  
-- Description:   
-- 
-- VHDL Test Bench Created by ISE for module: UARTtop
-- 
-- Dependencies:
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
--
-- Notes: 
-- This testbench has been automatically generated using types std_logic and
-- std_logic_vector for the ports of the unit under test.  Xilinx recommends
-- that these types always be used for the top-level I/O of a design in order
-- to guarantee that the testbench will bind correctly to the post-implementation 
-- simulation model.
--------------------------------------------------------------------------------
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
 
-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--USE ieee.numeric_std.ALL;
 
ENTITY UARTtb IS
END UARTtb;
 
ARCHITECTURE behavior OF UARTtb IS 
 
    -- Component Declaration for the Unit Under Test (UUT)
 
    COMPONENT UARTtop
    PORT(
         clk : IN  std_logic;
         reset : IN  std_logic;
         rx : IN  std_logic;
         tx : OUT  std_logic
        );
    END COMPONENT;
    

   --Inputs
   signal clk : std_logic := '0';
   signal reset : std_logic := '0';
   signal rx : std_logic := '1';

 	--Outputs
   signal tx : std_logic;

   -- Clock period definitions
   constant clk_period : time := 0.000037 ms;
 
BEGIN
 
	-- Instantiate the Unit Under Test (UUT)
   uut: UARTtop PORT MAP (
          clk => clk,
          reset => reset,
          rx => rx,
          tx => tx
        );

   -- Clock process definitions
   clk_process :process
   begin
		clk <= '0';
		wait for clk_period/2;
		clk <= '1';
		wait for clk_period/2;
   end process;
 

   -- Stimulus process
   stim_proc: process
   begin		
      -- hold reset state for 100 ns.
      wait for 100 ns;	
		
		rx <='0';		--start
      wait for 103600 ns;
		rx <= '1';		--prvi bit
		wait for 103600 ns;
		rx <= '0';
		wait for 103600 ns;
		rx <= '0';
		wait for 103600 ns;
		rx <= '0';
		wait for 103600 ns;
		rx <= '1';
		wait for 103600 ns;
		rx <= '1';
		wait for 103600 ns;
		rx <= '0';
		wait for 103600 ns;
		rx <= '0';		--zadnji
		wait for 103600 ns;
		rx <= '1';			-- stop
		
		wait for 103600 ns;
		rx <='0';			--start
      wait for 103600 ns;
		rx <= '1';			--prvi bit
		wait for 103600 ns;
		rx <= '1';
		wait for 103600 ns;
		rx <= '0';
		wait for 103600 ns;
		rx <= '0';
		wait for 103600 ns;
		rx <= '1';
		wait for 103600 ns;
		rx <= '0';
		wait for 103600 ns;
		rx <= '0';
		wait for 103600 ns;
		rx <= '0';		--zadnji
		wait for 103600 ns;
		rx <= '1';		-- stop
      -- insert stimulus here 

      wait;
   end process;

END;
